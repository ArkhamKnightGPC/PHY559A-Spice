.include cmosws.mod
			
Vsd 2 0 dc 3.3V
Vsg 2 1 dc 1V
M1  0 1 2 2 MODP L=0.6U W=6.0U
			
.dc Vsd 0 3.3 50mV Vsg 1 3 1V
.end