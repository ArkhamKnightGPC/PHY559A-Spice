.include cmosws.mod
			
Vdd 1 0 dc 3.3V
Va  2 0 dc 3.3V
Vb  3 0 dc 1.0V
M1  1 2 4 1 MODP L=0.6U W=6.0U
M2  1 3 4 1 MODP L=0.6U W=6.0U
M3  4 2 5 0 MODN L=0.6U W=6.0U
M4  5 3 0 0 MODN L=0.6U W=6.0U
			
.dc Vb 0 3.3 50mV
.end