.include cmosws.mod
*.include cmostm.mod

.option temp = -40
*.option temp = 125

Vin 1 0 pulse(0.0V 3.3V 5ns 1ns 1ns 3ns 8ns)
Vdd 2 0 dc 3.3V
M1  3 1 0 0 MODN L=0.6U W=3.0U
M2  2 1 3 2 MODP L=0.6U W=6.0U
C1  3 0 0.5pF

.tran 0.05ns 16ns
.end