.include cmosws.mod
			
Vin 1 0 dc 1V
Vdd 2 0 dc 3.3V
M1  3 1 0 0 MODN L=0.6U W=3.0U
M2  2 1 3 2 MODP L=0.6U W=12.0U
	
.dc Vin 0 3.3 50mV
.end